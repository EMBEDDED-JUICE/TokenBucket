/* Write a Verilog module named token_bucket that implements a token bucket rate limiter.
Parameters:

DEN (default 16): denominator for fractional rate control (tokens per request).

RATE_NUM (default 3): number of tokens added per cycle.

BURST_MAX (default 8): maximum burst size, expressed in requests.

TOKEN_COST (default = DEN): tokens consumed per granted request.

Inputs:

clk: clock.

rst_n: active-low synchronous reset.

req_i: request input.

Outputs:

grant_o: asserted when a request is accepted and tokens are consumed.

ready_o: asserted whenever enough tokens are available for a request.

Functional Behavior:

Maintain an internal token counter (width at least 32 bits).

On every clock cycle, add RATE_NUM tokens, but do not exceed the maximum capacity (BURST_MAX * DEN).

If req_i is high and tokens ≥ TOKEN_COST:

Assert grant_o for one cycle.

Subtract TOKEN_COST tokens.

Otherwise, keep grant_o low.

ready_o is high whenever tokens ≥ TOKEN_COST.

On reset (rst_n = 0), initialize the token counter to full capacity (BURST_MAX * DEN) and clear grant_o.*/

module top_module #(
    parameter DEN = 16,
    parameter RATE_NUM = 3,
    parameter BURST_MAX = 8,
    parameter TOKEN_COST = DEN
) (
    input  wire clk,
    input  wire rst_n,
    input  wire req_i,
    output wire grant_o,
    output wire ready_o
);

    // Implement the token bucket as specified above.

endmodule
